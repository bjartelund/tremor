﻿Movement,Anomaly
10089,0
10107,0
10086,0
10099,0
12417,1
10095,0
11009,1
12225,1
10158,0
16741,1
22189,1
19938,1
21431,1
9846,0
10211,0
10266,0
11884,1
12659,1
10433,0
19668,1
15896,1
11310,1
16359,1
